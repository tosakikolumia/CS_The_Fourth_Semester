`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/04/02 12:31:28
// Design Name: 
// Module Name: MULTU_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MULTU_tb;
    reg [31:0] a, b;
    wire [63:0] product;
    reg clk;
    reg reset;
    // 实例化 MULTU 模块
    MULTU uut (
        .clk(clk), // 时钟信号
        .reset(reset), // 复位信号
        .a(a),
        .b(b),
        .z(product)
    );
    
    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // 复位信号置位
        reset = 1'b1;
        #10;
        reset = 1'b0;
        #10;
        a = 32'b11111111111111111111111111111111; b = 32'b11111111111111111111111111111111;
        #10;
        // 测试用例
        a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000000;
        #10;
        a = 32'b00000000000000000000000010110011; b = 32'b00000000000000000000000000000000;
        #10;
        a = 32'b00000000000000000000000011111111; b = 32'b00000000000000000000000011111111;
        #10;
        a = 32'b00000000000000000000000010000000; b = 32'b00000000000000000000000010101010;
        #10;
        a = 32'b00000000000000000000000010101010; b = 32'b00000000000000000000000010000000;
        #10;
        a = 32'b00000000000000000000000000101101; b = 32'b00000000000000000000000011010000;
        #10;
        a = 32'b0000000000000000000000001000111; b = 32'b00000000000000000000000000001110;
        #10;
        
    end

endmodule
