`timescale 1ns / 1ps  
module MULT_tb;  
    reg clk; // 乘法器时钟信号  
    reg reset; // 复位信号，高电平有效  
    reg [31:0] a; // 输入 a (被乘数)  
    reg [31:0] b; // 输入 b (乘数)  
    wire [63:0] z; // 乘积输出 z  

    initial begin  
        clk = 0;  
        forever #10 clk = ~clk; 
    end  

    initial begin  
        reset = 1;  
        #100;  
        reset = 0;  
        a = 0;  
        b = 0;  
        
        #100;  
        a = 0;   
        b = 32'b1111_1111_1111_1111_1111_1111_1111_1111; // Test case 1  
        #100;  
        
        a = 32'b1000_0000_0000_0000_0000_0000_1011_0011; // Test case 2  
        b = 0;  
        #100;  
        
        a = 32'b1111_1111_1111_1111_1111_1111_1111_1111; // Test case 3  
        b = 32'b1111_1111_1111_1111_1111_1111_1111_1111;  
        #100;  
        
        a = 32'b1000_0000_0000_0000_0000_0000_1000_0000; // Test case 4  
        b = 32'b0000_0000_0000_0000_0000_0000_1010_1010;  
        #100;  
        
        a = 32'b0000_0000_0000_0000_0000_0000_1010_1010; // Test case 5  
        b = 32'b1000_0000_0000_0000_0000_0000_1000_0000;  
        #100;  
        
        a = 32'b0000_0000_0000_0000_0000_0000_1110_1101; // Test case 6  
        b = 32'b0000_0000_0000_0000_0000_0000_1101_0000;  
        #100;  
        
        a = 32'b0000_0000_0000_0000_0000_0000_1000_1111; // Test case 7  
        b = 32'b0000_0000_0000_0000_0000_0000_0000_1110;  
    end  

    MULT 
    MULT_init(  
        .clk(clk),  
        .reset(reset),  
        .a(a),  
        .b(b),  
        .z(z)  
    );  
endmodule  